-- qsys.vhd

-- Generated using ACDS version 20.1 720

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity qsys is
	port (
		btn_export    : in    std_logic_vector(7 downto 0)  := (others => '0'); --     btn.export
		clk_clk       : in    std_logic                     := '0';             --     clk.clk
		d7seg_export  : out   std_logic_vector(15 downto 0);                    --   d7seg.export
		eeprom_sda_in : in    std_logic                     := '0';             --  eeprom.sda_in
		eeprom_scl_in : in    std_logic                     := '0';             --        .scl_in
		eeprom_sda_oe : out   std_logic;                                        --        .sda_oe
		eeprom_scl_oe : out   std_logic;                                        --        .scl_oe
		enc_spi_MISO  : in    std_logic                     := '0';             -- enc_spi.MISO
		enc_spi_MOSI  : out   std_logic;                                        --        .MOSI
		enc_spi_SCLK  : out   std_logic;                                        --        .SCLK
		enc_spi_SS_n  : out   std_logic;                                        --        .SS_n
		led_export    : out   std_logic_vector(3 downto 0);                     --     led.export
		ram_addr      : out   std_logic_vector(11 downto 0);                    --     ram.addr
		ram_ba        : out   std_logic_vector(1 downto 0);                     --        .ba
		ram_cas_n     : out   std_logic;                                        --        .cas_n
		ram_cke       : out   std_logic;                                        --        .cke
		ram_cs_n      : out   std_logic;                                        --        .cs_n
		ram_dq        : inout std_logic_vector(15 downto 0) := (others => '0'); --        .dq
		ram_dqm       : out   std_logic_vector(1 downto 0);                     --        .dqm
		ram_ras_n     : out   std_logic;                                        --        .ras_n
		ram_we_n      : out   std_logic;                                        --        .we_n
		reset_reset_n : in    std_logic                     := '0';             --   reset.reset_n
		temp_sda_in   : in    std_logic                     := '0';             --    temp.sda_in
		temp_scl_in   : in    std_logic                     := '0';             --        .scl_in
		temp_sda_oe   : out   std_logic;                                        --        .sda_oe
		temp_scl_oe   : out   std_logic                                         --        .scl_oe
	);
end entity qsys;

architecture rtl of qsys is
	component altera_avalon_i2c is
		generic (
			USE_AV_ST       : integer := 0;
			FIFO_DEPTH      : integer := 4;
			FIFO_DEPTH_LOG2 : integer := 2
		);
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			rst_n     : in  std_logic                     := 'X';             -- reset_n
			intr      : out std_logic;                                        -- irq
			addr      : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			sda_in    : in  std_logic                     := 'X';             -- sda_in
			scl_in    : in  std_logic                     := 'X';             -- scl_in
			sda_oe    : out std_logic;                                        -- sda_oe
			scl_oe    : out std_logic;                                        -- scl_oe
			src_data  : out std_logic_vector(7 downto 0);                     -- data
			src_valid : out std_logic;                                        -- valid
			src_ready : in  std_logic                     := 'X';             -- ready
			snk_data  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data
			snk_valid : in  std_logic                     := 'X';             -- valid
			snk_ready : out std_logic                                         -- ready
		);
	end component altera_avalon_i2c;

	component qsys_JTAG_UART is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component qsys_JTAG_UART;

	component qsys_NIOSII is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(24 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(24 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component qsys_NIOSII;

	component qsys_PIO_BTN is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component qsys_PIO_BTN;

	component qsys_PIO_D7SEG is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component qsys_PIO_D7SEG;

	component qsys_PIO_LED is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(3 downto 0)                      -- export
		);
	end component qsys_PIO_LED;

	component qsys_RAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(21 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(11 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component qsys_RAM;

	component qsys_SPI_MASTER is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component qsys_SPI_MASTER;

	component qsys_SYSID is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component qsys_SYSID;

	component qsys_SYS_TIMER is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component qsys_SYS_TIMER;

	component qsys_TS_TIMER is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component qsys_TS_TIMER;

	component qsys_mm_interconnect_0 is
		port (
			clk_0_clk_clk                            : in  std_logic                     := 'X';             -- clk
			NIOSII_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			NIOSII_data_master_address               : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			NIOSII_data_master_waitrequest           : out std_logic;                                        -- waitrequest
			NIOSII_data_master_byteenable            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			NIOSII_data_master_read                  : in  std_logic                     := 'X';             -- read
			NIOSII_data_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			NIOSII_data_master_write                 : in  std_logic                     := 'X';             -- write
			NIOSII_data_master_writedata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			NIOSII_data_master_debugaccess           : in  std_logic                     := 'X';             -- debugaccess
			NIOSII_instruction_master_address        : in  std_logic_vector(24 downto 0) := (others => 'X'); -- address
			NIOSII_instruction_master_waitrequest    : out std_logic;                                        -- waitrequest
			NIOSII_instruction_master_read           : in  std_logic                     := 'X';             -- read
			NIOSII_instruction_master_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			I2C_EEPROM_csr_address                   : out std_logic_vector(3 downto 0);                     -- address
			I2C_EEPROM_csr_write                     : out std_logic;                                        -- write
			I2C_EEPROM_csr_read                      : out std_logic;                                        -- read
			I2C_EEPROM_csr_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			I2C_EEPROM_csr_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			I2C_TEMP_csr_address                     : out std_logic_vector(3 downto 0);                     -- address
			I2C_TEMP_csr_write                       : out std_logic;                                        -- write
			I2C_TEMP_csr_read                        : out std_logic;                                        -- read
			I2C_TEMP_csr_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			I2C_TEMP_csr_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_address      : out std_logic_vector(0 downto 0);                     -- address
			JTAG_UART_avalon_jtag_slave_write        : out std_logic;                                        -- write
			JTAG_UART_avalon_jtag_slave_read         : out std_logic;                                        -- read
			JTAG_UART_avalon_jtag_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_UART_avalon_jtag_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_UART_avalon_jtag_slave_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect   : out std_logic;                                        -- chipselect
			NIOSII_debug_mem_slave_address           : out std_logic_vector(8 downto 0);                     -- address
			NIOSII_debug_mem_slave_write             : out std_logic;                                        -- write
			NIOSII_debug_mem_slave_read              : out std_logic;                                        -- read
			NIOSII_debug_mem_slave_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			NIOSII_debug_mem_slave_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			NIOSII_debug_mem_slave_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			NIOSII_debug_mem_slave_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			NIOSII_debug_mem_slave_debugaccess       : out std_logic;                                        -- debugaccess
			PIO_BTN_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			PIO_BTN_s1_write                         : out std_logic;                                        -- write
			PIO_BTN_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIO_BTN_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			PIO_BTN_s1_chipselect                    : out std_logic;                                        -- chipselect
			PIO_D7SEG_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			PIO_D7SEG_s1_write                       : out std_logic;                                        -- write
			PIO_D7SEG_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIO_D7SEG_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			PIO_D7SEG_s1_chipselect                  : out std_logic;                                        -- chipselect
			PIO_LED_s1_address                       : out std_logic_vector(1 downto 0);                     -- address
			PIO_LED_s1_write                         : out std_logic;                                        -- write
			PIO_LED_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PIO_LED_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			PIO_LED_s1_chipselect                    : out std_logic;                                        -- chipselect
			RAM_s1_address                           : out std_logic_vector(21 downto 0);                    -- address
			RAM_s1_write                             : out std_logic;                                        -- write
			RAM_s1_read                              : out std_logic;                                        -- read
			RAM_s1_readdata                          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			RAM_s1_writedata                         : out std_logic_vector(15 downto 0);                    -- writedata
			RAM_s1_byteenable                        : out std_logic_vector(1 downto 0);                     -- byteenable
			RAM_s1_readdatavalid                     : in  std_logic                     := 'X';             -- readdatavalid
			RAM_s1_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			RAM_s1_chipselect                        : out std_logic;                                        -- chipselect
			SPI_MASTER_spi_control_port_address      : out std_logic_vector(2 downto 0);                     -- address
			SPI_MASTER_spi_control_port_write        : out std_logic;                                        -- write
			SPI_MASTER_spi_control_port_read         : out std_logic;                                        -- read
			SPI_MASTER_spi_control_port_readdata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SPI_MASTER_spi_control_port_writedata    : out std_logic_vector(15 downto 0);                    -- writedata
			SPI_MASTER_spi_control_port_chipselect   : out std_logic;                                        -- chipselect
			SYS_TIMER_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			SYS_TIMER_s1_write                       : out std_logic;                                        -- write
			SYS_TIMER_s1_readdata                    : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SYS_TIMER_s1_writedata                   : out std_logic_vector(15 downto 0);                    -- writedata
			SYS_TIMER_s1_chipselect                  : out std_logic;                                        -- chipselect
			SYSID_control_slave_address              : out std_logic_vector(0 downto 0);                     -- address
			SYSID_control_slave_readdata             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TS_TIMER_s1_address                      : out std_logic_vector(2 downto 0);                     -- address
			TS_TIMER_s1_write                        : out std_logic;                                        -- write
			TS_TIMER_s1_readdata                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			TS_TIMER_s1_writedata                    : out std_logic_vector(15 downto 0);                    -- writedata
			TS_TIMER_s1_chipselect                   : out std_logic                                         -- chipselect
		);
	end component qsys_mm_interconnect_0;

	component qsys_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component qsys_irq_mapper;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal niosii_data_master_readdata                                   : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOSII_data_master_readdata -> NIOSII:d_readdata
	signal niosii_data_master_waitrequest                                : std_logic;                     -- mm_interconnect_0:NIOSII_data_master_waitrequest -> NIOSII:d_waitrequest
	signal niosii_data_master_debugaccess                                : std_logic;                     -- NIOSII:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOSII_data_master_debugaccess
	signal niosii_data_master_address                                    : std_logic_vector(24 downto 0); -- NIOSII:d_address -> mm_interconnect_0:NIOSII_data_master_address
	signal niosii_data_master_byteenable                                 : std_logic_vector(3 downto 0);  -- NIOSII:d_byteenable -> mm_interconnect_0:NIOSII_data_master_byteenable
	signal niosii_data_master_read                                       : std_logic;                     -- NIOSII:d_read -> mm_interconnect_0:NIOSII_data_master_read
	signal niosii_data_master_write                                      : std_logic;                     -- NIOSII:d_write -> mm_interconnect_0:NIOSII_data_master_write
	signal niosii_data_master_writedata                                  : std_logic_vector(31 downto 0); -- NIOSII:d_writedata -> mm_interconnect_0:NIOSII_data_master_writedata
	signal niosii_instruction_master_readdata                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOSII_instruction_master_readdata -> NIOSII:i_readdata
	signal niosii_instruction_master_waitrequest                         : std_logic;                     -- mm_interconnect_0:NIOSII_instruction_master_waitrequest -> NIOSII:i_waitrequest
	signal niosii_instruction_master_address                             : std_logic_vector(24 downto 0); -- NIOSII:i_address -> mm_interconnect_0:NIOSII_instruction_master_address
	signal niosii_instruction_master_read                                : std_logic;                     -- NIOSII:i_read -> mm_interconnect_0:NIOSII_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_chipselect -> JTAG_UART:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- JTAG_UART:av_readdata -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- JTAG_UART:av_waitrequest -> mm_interconnect_0:JTAG_UART_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_address -> JTAG_UART:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_UART_avalon_jtag_slave_writedata -> JTAG_UART:av_writedata
	signal mm_interconnect_0_sysid_control_slave_readdata                : std_logic_vector(31 downto 0); -- SYSID:readdata -> mm_interconnect_0:SYSID_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:SYSID_control_slave_address -> SYSID:address
	signal mm_interconnect_0_i2c_temp_csr_readdata                       : std_logic_vector(31 downto 0); -- I2C_TEMP:readdata -> mm_interconnect_0:I2C_TEMP_csr_readdata
	signal mm_interconnect_0_i2c_temp_csr_address                        : std_logic_vector(3 downto 0);  -- mm_interconnect_0:I2C_TEMP_csr_address -> I2C_TEMP:addr
	signal mm_interconnect_0_i2c_temp_csr_read                           : std_logic;                     -- mm_interconnect_0:I2C_TEMP_csr_read -> I2C_TEMP:read
	signal mm_interconnect_0_i2c_temp_csr_write                          : std_logic;                     -- mm_interconnect_0:I2C_TEMP_csr_write -> I2C_TEMP:write
	signal mm_interconnect_0_i2c_temp_csr_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:I2C_TEMP_csr_writedata -> I2C_TEMP:writedata
	signal mm_interconnect_0_i2c_eeprom_csr_readdata                     : std_logic_vector(31 downto 0); -- I2C_EEPROM:readdata -> mm_interconnect_0:I2C_EEPROM_csr_readdata
	signal mm_interconnect_0_i2c_eeprom_csr_address                      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:I2C_EEPROM_csr_address -> I2C_EEPROM:addr
	signal mm_interconnect_0_i2c_eeprom_csr_read                         : std_logic;                     -- mm_interconnect_0:I2C_EEPROM_csr_read -> I2C_EEPROM:read
	signal mm_interconnect_0_i2c_eeprom_csr_write                        : std_logic;                     -- mm_interconnect_0:I2C_EEPROM_csr_write -> I2C_EEPROM:write
	signal mm_interconnect_0_i2c_eeprom_csr_writedata                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:I2C_EEPROM_csr_writedata -> I2C_EEPROM:writedata
	signal mm_interconnect_0_niosii_debug_mem_slave_readdata             : std_logic_vector(31 downto 0); -- NIOSII:debug_mem_slave_readdata -> mm_interconnect_0:NIOSII_debug_mem_slave_readdata
	signal mm_interconnect_0_niosii_debug_mem_slave_waitrequest          : std_logic;                     -- NIOSII:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOSII_debug_mem_slave_waitrequest
	signal mm_interconnect_0_niosii_debug_mem_slave_debugaccess          : std_logic;                     -- mm_interconnect_0:NIOSII_debug_mem_slave_debugaccess -> NIOSII:debug_mem_slave_debugaccess
	signal mm_interconnect_0_niosii_debug_mem_slave_address              : std_logic_vector(8 downto 0);  -- mm_interconnect_0:NIOSII_debug_mem_slave_address -> NIOSII:debug_mem_slave_address
	signal mm_interconnect_0_niosii_debug_mem_slave_read                 : std_logic;                     -- mm_interconnect_0:NIOSII_debug_mem_slave_read -> NIOSII:debug_mem_slave_read
	signal mm_interconnect_0_niosii_debug_mem_slave_byteenable           : std_logic_vector(3 downto 0);  -- mm_interconnect_0:NIOSII_debug_mem_slave_byteenable -> NIOSII:debug_mem_slave_byteenable
	signal mm_interconnect_0_niosii_debug_mem_slave_write                : std_logic;                     -- mm_interconnect_0:NIOSII_debug_mem_slave_write -> NIOSII:debug_mem_slave_write
	signal mm_interconnect_0_niosii_debug_mem_slave_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:NIOSII_debug_mem_slave_writedata -> NIOSII:debug_mem_slave_writedata
	signal mm_interconnect_0_ram_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:RAM_s1_chipselect -> RAM:az_cs
	signal mm_interconnect_0_ram_s1_readdata                             : std_logic_vector(15 downto 0); -- RAM:za_data -> mm_interconnect_0:RAM_s1_readdata
	signal mm_interconnect_0_ram_s1_waitrequest                          : std_logic;                     -- RAM:za_waitrequest -> mm_interconnect_0:RAM_s1_waitrequest
	signal mm_interconnect_0_ram_s1_address                              : std_logic_vector(21 downto 0); -- mm_interconnect_0:RAM_s1_address -> RAM:az_addr
	signal mm_interconnect_0_ram_s1_read                                 : std_logic;                     -- mm_interconnect_0:RAM_s1_read -> mm_interconnect_0_ram_s1_read:in
	signal mm_interconnect_0_ram_s1_byteenable                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:RAM_s1_byteenable -> mm_interconnect_0_ram_s1_byteenable:in
	signal mm_interconnect_0_ram_s1_readdatavalid                        : std_logic;                     -- RAM:za_valid -> mm_interconnect_0:RAM_s1_readdatavalid
	signal mm_interconnect_0_ram_s1_write                                : std_logic;                     -- mm_interconnect_0:RAM_s1_write -> mm_interconnect_0_ram_s1_write:in
	signal mm_interconnect_0_ram_s1_writedata                            : std_logic_vector(15 downto 0); -- mm_interconnect_0:RAM_s1_writedata -> RAM:az_data
	signal mm_interconnect_0_pio_led_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:PIO_LED_s1_chipselect -> PIO_LED:chipselect
	signal mm_interconnect_0_pio_led_s1_readdata                         : std_logic_vector(31 downto 0); -- PIO_LED:readdata -> mm_interconnect_0:PIO_LED_s1_readdata
	signal mm_interconnect_0_pio_led_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIO_LED_s1_address -> PIO_LED:address
	signal mm_interconnect_0_pio_led_s1_write                            : std_logic;                     -- mm_interconnect_0:PIO_LED_s1_write -> mm_interconnect_0_pio_led_s1_write:in
	signal mm_interconnect_0_pio_led_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:PIO_LED_s1_writedata -> PIO_LED:writedata
	signal mm_interconnect_0_pio_btn_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:PIO_BTN_s1_chipselect -> PIO_BTN:chipselect
	signal mm_interconnect_0_pio_btn_s1_readdata                         : std_logic_vector(31 downto 0); -- PIO_BTN:readdata -> mm_interconnect_0:PIO_BTN_s1_readdata
	signal mm_interconnect_0_pio_btn_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIO_BTN_s1_address -> PIO_BTN:address
	signal mm_interconnect_0_pio_btn_s1_write                            : std_logic;                     -- mm_interconnect_0:PIO_BTN_s1_write -> mm_interconnect_0_pio_btn_s1_write:in
	signal mm_interconnect_0_pio_btn_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:PIO_BTN_s1_writedata -> PIO_BTN:writedata
	signal mm_interconnect_0_sys_timer_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:SYS_TIMER_s1_chipselect -> SYS_TIMER:chipselect
	signal mm_interconnect_0_sys_timer_s1_readdata                       : std_logic_vector(15 downto 0); -- SYS_TIMER:readdata -> mm_interconnect_0:SYS_TIMER_s1_readdata
	signal mm_interconnect_0_sys_timer_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SYS_TIMER_s1_address -> SYS_TIMER:address
	signal mm_interconnect_0_sys_timer_s1_write                          : std_logic;                     -- mm_interconnect_0:SYS_TIMER_s1_write -> mm_interconnect_0_sys_timer_s1_write:in
	signal mm_interconnect_0_sys_timer_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:SYS_TIMER_s1_writedata -> SYS_TIMER:writedata
	signal mm_interconnect_0_ts_timer_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:TS_TIMER_s1_chipselect -> TS_TIMER:chipselect
	signal mm_interconnect_0_ts_timer_s1_readdata                        : std_logic_vector(15 downto 0); -- TS_TIMER:readdata -> mm_interconnect_0:TS_TIMER_s1_readdata
	signal mm_interconnect_0_ts_timer_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:TS_TIMER_s1_address -> TS_TIMER:address
	signal mm_interconnect_0_ts_timer_s1_write                           : std_logic;                     -- mm_interconnect_0:TS_TIMER_s1_write -> mm_interconnect_0_ts_timer_s1_write:in
	signal mm_interconnect_0_ts_timer_s1_writedata                       : std_logic_vector(15 downto 0); -- mm_interconnect_0:TS_TIMER_s1_writedata -> TS_TIMER:writedata
	signal mm_interconnect_0_pio_d7seg_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:PIO_D7SEG_s1_chipselect -> PIO_D7SEG:chipselect
	signal mm_interconnect_0_pio_d7seg_s1_readdata                       : std_logic_vector(31 downto 0); -- PIO_D7SEG:readdata -> mm_interconnect_0:PIO_D7SEG_s1_readdata
	signal mm_interconnect_0_pio_d7seg_s1_address                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PIO_D7SEG_s1_address -> PIO_D7SEG:address
	signal mm_interconnect_0_pio_d7seg_s1_write                          : std_logic;                     -- mm_interconnect_0:PIO_D7SEG_s1_write -> mm_interconnect_0_pio_d7seg_s1_write:in
	signal mm_interconnect_0_pio_d7seg_s1_writedata                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:PIO_D7SEG_s1_writedata -> PIO_D7SEG:writedata
	signal mm_interconnect_0_spi_master_spi_control_port_chipselect      : std_logic;                     -- mm_interconnect_0:SPI_MASTER_spi_control_port_chipselect -> SPI_MASTER:spi_select
	signal mm_interconnect_0_spi_master_spi_control_port_readdata        : std_logic_vector(15 downto 0); -- SPI_MASTER:data_to_cpu -> mm_interconnect_0:SPI_MASTER_spi_control_port_readdata
	signal mm_interconnect_0_spi_master_spi_control_port_address         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:SPI_MASTER_spi_control_port_address -> SPI_MASTER:mem_addr
	signal mm_interconnect_0_spi_master_spi_control_port_read            : std_logic;                     -- mm_interconnect_0:SPI_MASTER_spi_control_port_read -> mm_interconnect_0_spi_master_spi_control_port_read:in
	signal mm_interconnect_0_spi_master_spi_control_port_write           : std_logic;                     -- mm_interconnect_0:SPI_MASTER_spi_control_port_write -> mm_interconnect_0_spi_master_spi_control_port_write:in
	signal mm_interconnect_0_spi_master_spi_control_port_writedata       : std_logic_vector(15 downto 0); -- mm_interconnect_0:SPI_MASTER_spi_control_port_writedata -> SPI_MASTER:data_from_cpu
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- SYS_TIMER:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- JTAG_UART:av_irq -> irq_mapper:receiver1_irq
	signal niosii_irq_irq                                                : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> NIOSII:irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:NIOSII_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [NIOSII:reset_req, rst_translator:reset_req_in]
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> rst_controller:reset_in0
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> JTAG_UART:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> JTAG_UART:av_write_n
	signal mm_interconnect_0_ram_s1_read_ports_inv                       : std_logic;                     -- mm_interconnect_0_ram_s1_read:inv -> RAM:az_rd_n
	signal mm_interconnect_0_ram_s1_byteenable_ports_inv                 : std_logic_vector(1 downto 0);  -- mm_interconnect_0_ram_s1_byteenable:inv -> RAM:az_be_n
	signal mm_interconnect_0_ram_s1_write_ports_inv                      : std_logic;                     -- mm_interconnect_0_ram_s1_write:inv -> RAM:az_wr_n
	signal mm_interconnect_0_pio_led_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_pio_led_s1_write:inv -> PIO_LED:write_n
	signal mm_interconnect_0_pio_btn_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_pio_btn_s1_write:inv -> PIO_BTN:write_n
	signal mm_interconnect_0_sys_timer_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_sys_timer_s1_write:inv -> SYS_TIMER:write_n
	signal mm_interconnect_0_ts_timer_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_ts_timer_s1_write:inv -> TS_TIMER:write_n
	signal mm_interconnect_0_pio_d7seg_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_pio_d7seg_s1_write:inv -> PIO_D7SEG:write_n
	signal mm_interconnect_0_spi_master_spi_control_port_read_ports_inv  : std_logic;                     -- mm_interconnect_0_spi_master_spi_control_port_read:inv -> SPI_MASTER:read_n
	signal mm_interconnect_0_spi_master_spi_control_port_write_ports_inv : std_logic;                     -- mm_interconnect_0_spi_master_spi_control_port_write:inv -> SPI_MASTER:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [I2C_EEPROM:rst_n, I2C_TEMP:rst_n, JTAG_UART:rst_n, NIOSII:reset_n, PIO_BTN:reset_n, PIO_D7SEG:reset_n, PIO_LED:reset_n, RAM:reset_n, SPI_MASTER:reset_n, SYSID:reset_n, SYS_TIMER:reset_n, TS_TIMER:reset_n]

begin

	i2c_eeprom : component altera_avalon_i2c
		generic map (
			USE_AV_ST       => 0,
			FIFO_DEPTH      => 8,
			FIFO_DEPTH_LOG2 => 3
		)
		port map (
			clk       => clk_clk,                                    --            clock.clk
			rst_n     => rst_controller_reset_out_reset_ports_inv,   --       reset_sink.reset_n
			intr      => open,                                       -- interrupt_sender.irq
			addr      => mm_interconnect_0_i2c_eeprom_csr_address,   --              csr.address
			read      => mm_interconnect_0_i2c_eeprom_csr_read,      --                 .read
			write     => mm_interconnect_0_i2c_eeprom_csr_write,     --                 .write
			writedata => mm_interconnect_0_i2c_eeprom_csr_writedata, --                 .writedata
			readdata  => mm_interconnect_0_i2c_eeprom_csr_readdata,  --                 .readdata
			sda_in    => eeprom_sda_in,                              --       i2c_serial.sda_in
			scl_in    => eeprom_scl_in,                              --                 .scl_in
			sda_oe    => eeprom_sda_oe,                              --                 .sda_oe
			scl_oe    => eeprom_scl_oe,                              --                 .scl_oe
			src_data  => open,                                       --      (terminated)
			src_valid => open,                                       --      (terminated)
			src_ready => '0',                                        --      (terminated)
			snk_data  => "0000000000000000",                         --      (terminated)
			snk_valid => '0',                                        --      (terminated)
			snk_ready => open                                        --      (terminated)
		);

	i2c_temp : component altera_avalon_i2c
		generic map (
			USE_AV_ST       => 0,
			FIFO_DEPTH      => 8,
			FIFO_DEPTH_LOG2 => 3
		)
		port map (
			clk       => clk_clk,                                  --            clock.clk
			rst_n     => rst_controller_reset_out_reset_ports_inv, --       reset_sink.reset_n
			intr      => open,                                     -- interrupt_sender.irq
			addr      => mm_interconnect_0_i2c_temp_csr_address,   --              csr.address
			read      => mm_interconnect_0_i2c_temp_csr_read,      --                 .read
			write     => mm_interconnect_0_i2c_temp_csr_write,     --                 .write
			writedata => mm_interconnect_0_i2c_temp_csr_writedata, --                 .writedata
			readdata  => mm_interconnect_0_i2c_temp_csr_readdata,  --                 .readdata
			sda_in    => temp_sda_in,                              --       i2c_serial.sda_in
			scl_in    => temp_scl_in,                              --                 .scl_in
			sda_oe    => temp_sda_oe,                              --                 .sda_oe
			scl_oe    => temp_scl_oe,                              --                 .scl_oe
			src_data  => open,                                     --      (terminated)
			src_valid => open,                                     --      (terminated)
			src_ready => '0',                                      --      (terminated)
			snk_data  => "0000000000000000",                       --      (terminated)
			snk_valid => '0',                                      --      (terminated)
			snk_ready => open                                      --      (terminated)
		);

	jtag_uart : component qsys_JTAG_UART
		port map (
			clk            => clk_clk,                                                       --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	niosii : component qsys_NIOSII
		port map (
			clk                                 => clk_clk,                                              --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,             --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                   --                          .reset_req
			d_address                           => niosii_data_master_address,                           --               data_master.address
			d_byteenable                        => niosii_data_master_byteenable,                        --                          .byteenable
			d_read                              => niosii_data_master_read,                              --                          .read
			d_readdata                          => niosii_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => niosii_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => niosii_data_master_write,                             --                          .write
			d_writedata                         => niosii_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => niosii_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => niosii_instruction_master_address,                    --        instruction_master.address
			i_read                              => niosii_instruction_master_read,                       --                          .read
			i_readdata                          => niosii_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => niosii_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => niosii_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => open,                                                 --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_niosii_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_niosii_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_niosii_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_niosii_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_niosii_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_niosii_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_niosii_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_niosii_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                  -- custom_instruction_master.readra
		);

	pio_btn : component qsys_PIO_BTN
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_btn_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_btn_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_btn_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_btn_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_btn_s1_readdata,        --                    .readdata
			in_port    => btn_export,                                   -- external_connection.export
			irq        => open                                          --                 irq.irq
		);

	pio_d7seg : component qsys_PIO_D7SEG
		port map (
			clk        => clk_clk,                                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       --               reset.reset_n
			address    => mm_interconnect_0_pio_d7seg_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_d7seg_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_d7seg_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_d7seg_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_d7seg_s1_readdata,        --                    .readdata
			out_port   => d7seg_export                                    -- external_connection.export
		);

	pio_led : component qsys_PIO_LED
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_led_s1_readdata,        --                    .readdata
			out_port   => led_export                                    -- external_connection.export
		);

	ram : component qsys_RAM
		port map (
			clk            => clk_clk,                                       --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,      -- reset.reset_n
			az_addr        => mm_interconnect_0_ram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_ram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_ram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_ram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_ram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_ram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_ram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_ram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_ram_s1_waitrequest,          --      .waitrequest
			zs_addr        => ram_addr,                                      --  wire.export
			zs_ba          => ram_ba,                                        --      .export
			zs_cas_n       => ram_cas_n,                                     --      .export
			zs_cke         => ram_cke,                                       --      .export
			zs_cs_n        => ram_cs_n,                                      --      .export
			zs_dq          => ram_dq,                                        --      .export
			zs_dqm         => ram_dqm,                                       --      .export
			zs_ras_n       => ram_ras_n,                                     --      .export
			zs_we_n        => ram_we_n                                       --      .export
		);

	spi_master : component qsys_SPI_MASTER
		port map (
			clk           => clk_clk,                                                       --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                      --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_master_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_master_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_master_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_master_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_master_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_master_spi_control_port_write_ports_inv, --                 .write_n
			irq           => open,                                                          --              irq.irq
			MISO          => enc_spi_MISO,                                                  --         external.export
			MOSI          => enc_spi_MOSI,                                                  --                 .export
			SCLK          => enc_spi_SCLK,                                                  --                 .export
			SS_n          => enc_spi_SS_n                                                   --                 .export
		);

	sysid : component qsys_SYSID
		port map (
			clock    => clk_clk,                                          --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	sys_timer : component qsys_SYS_TIMER
		port map (
			clk        => clk_clk,                                        --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       -- reset.reset_n
			address    => mm_interconnect_0_sys_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver0_irq                        --   irq.irq
		);

	ts_timer : component qsys_TS_TIMER
		port map (
			clk        => clk_clk,                                       --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      -- reset.reset_n
			address    => mm_interconnect_0_ts_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_ts_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_ts_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_ts_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_ts_timer_s1_write_ports_inv, --      .write_n
			irq        => open                                           --   irq.irq
		);

	mm_interconnect_0 : component qsys_mm_interconnect_0
		port map (
			clk_0_clk_clk                            => clk_clk,                                                   --                          clk_0_clk.clk
			NIOSII_reset_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- NIOSII_reset_reset_bridge_in_reset.reset
			NIOSII_data_master_address               => niosii_data_master_address,                                --                 NIOSII_data_master.address
			NIOSII_data_master_waitrequest           => niosii_data_master_waitrequest,                            --                                   .waitrequest
			NIOSII_data_master_byteenable            => niosii_data_master_byteenable,                             --                                   .byteenable
			NIOSII_data_master_read                  => niosii_data_master_read,                                   --                                   .read
			NIOSII_data_master_readdata              => niosii_data_master_readdata,                               --                                   .readdata
			NIOSII_data_master_write                 => niosii_data_master_write,                                  --                                   .write
			NIOSII_data_master_writedata             => niosii_data_master_writedata,                              --                                   .writedata
			NIOSII_data_master_debugaccess           => niosii_data_master_debugaccess,                            --                                   .debugaccess
			NIOSII_instruction_master_address        => niosii_instruction_master_address,                         --          NIOSII_instruction_master.address
			NIOSII_instruction_master_waitrequest    => niosii_instruction_master_waitrequest,                     --                                   .waitrequest
			NIOSII_instruction_master_read           => niosii_instruction_master_read,                            --                                   .read
			NIOSII_instruction_master_readdata       => niosii_instruction_master_readdata,                        --                                   .readdata
			I2C_EEPROM_csr_address                   => mm_interconnect_0_i2c_eeprom_csr_address,                  --                     I2C_EEPROM_csr.address
			I2C_EEPROM_csr_write                     => mm_interconnect_0_i2c_eeprom_csr_write,                    --                                   .write
			I2C_EEPROM_csr_read                      => mm_interconnect_0_i2c_eeprom_csr_read,                     --                                   .read
			I2C_EEPROM_csr_readdata                  => mm_interconnect_0_i2c_eeprom_csr_readdata,                 --                                   .readdata
			I2C_EEPROM_csr_writedata                 => mm_interconnect_0_i2c_eeprom_csr_writedata,                --                                   .writedata
			I2C_TEMP_csr_address                     => mm_interconnect_0_i2c_temp_csr_address,                    --                       I2C_TEMP_csr.address
			I2C_TEMP_csr_write                       => mm_interconnect_0_i2c_temp_csr_write,                      --                                   .write
			I2C_TEMP_csr_read                        => mm_interconnect_0_i2c_temp_csr_read,                       --                                   .read
			I2C_TEMP_csr_readdata                    => mm_interconnect_0_i2c_temp_csr_readdata,                   --                                   .readdata
			I2C_TEMP_csr_writedata                   => mm_interconnect_0_i2c_temp_csr_writedata,                  --                                   .writedata
			JTAG_UART_avalon_jtag_slave_address      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --        JTAG_UART_avalon_jtag_slave.address
			JTAG_UART_avalon_jtag_slave_write        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                   .write
			JTAG_UART_avalon_jtag_slave_read         => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                   .read
			JTAG_UART_avalon_jtag_slave_readdata     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                   .readdata
			JTAG_UART_avalon_jtag_slave_writedata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                   .writedata
			JTAG_UART_avalon_jtag_slave_waitrequest  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                   .waitrequest
			JTAG_UART_avalon_jtag_slave_chipselect   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                   .chipselect
			NIOSII_debug_mem_slave_address           => mm_interconnect_0_niosii_debug_mem_slave_address,          --             NIOSII_debug_mem_slave.address
			NIOSII_debug_mem_slave_write             => mm_interconnect_0_niosii_debug_mem_slave_write,            --                                   .write
			NIOSII_debug_mem_slave_read              => mm_interconnect_0_niosii_debug_mem_slave_read,             --                                   .read
			NIOSII_debug_mem_slave_readdata          => mm_interconnect_0_niosii_debug_mem_slave_readdata,         --                                   .readdata
			NIOSII_debug_mem_slave_writedata         => mm_interconnect_0_niosii_debug_mem_slave_writedata,        --                                   .writedata
			NIOSII_debug_mem_slave_byteenable        => mm_interconnect_0_niosii_debug_mem_slave_byteenable,       --                                   .byteenable
			NIOSII_debug_mem_slave_waitrequest       => mm_interconnect_0_niosii_debug_mem_slave_waitrequest,      --                                   .waitrequest
			NIOSII_debug_mem_slave_debugaccess       => mm_interconnect_0_niosii_debug_mem_slave_debugaccess,      --                                   .debugaccess
			PIO_BTN_s1_address                       => mm_interconnect_0_pio_btn_s1_address,                      --                         PIO_BTN_s1.address
			PIO_BTN_s1_write                         => mm_interconnect_0_pio_btn_s1_write,                        --                                   .write
			PIO_BTN_s1_readdata                      => mm_interconnect_0_pio_btn_s1_readdata,                     --                                   .readdata
			PIO_BTN_s1_writedata                     => mm_interconnect_0_pio_btn_s1_writedata,                    --                                   .writedata
			PIO_BTN_s1_chipselect                    => mm_interconnect_0_pio_btn_s1_chipselect,                   --                                   .chipselect
			PIO_D7SEG_s1_address                     => mm_interconnect_0_pio_d7seg_s1_address,                    --                       PIO_D7SEG_s1.address
			PIO_D7SEG_s1_write                       => mm_interconnect_0_pio_d7seg_s1_write,                      --                                   .write
			PIO_D7SEG_s1_readdata                    => mm_interconnect_0_pio_d7seg_s1_readdata,                   --                                   .readdata
			PIO_D7SEG_s1_writedata                   => mm_interconnect_0_pio_d7seg_s1_writedata,                  --                                   .writedata
			PIO_D7SEG_s1_chipselect                  => mm_interconnect_0_pio_d7seg_s1_chipselect,                 --                                   .chipselect
			PIO_LED_s1_address                       => mm_interconnect_0_pio_led_s1_address,                      --                         PIO_LED_s1.address
			PIO_LED_s1_write                         => mm_interconnect_0_pio_led_s1_write,                        --                                   .write
			PIO_LED_s1_readdata                      => mm_interconnect_0_pio_led_s1_readdata,                     --                                   .readdata
			PIO_LED_s1_writedata                     => mm_interconnect_0_pio_led_s1_writedata,                    --                                   .writedata
			PIO_LED_s1_chipselect                    => mm_interconnect_0_pio_led_s1_chipselect,                   --                                   .chipselect
			RAM_s1_address                           => mm_interconnect_0_ram_s1_address,                          --                             RAM_s1.address
			RAM_s1_write                             => mm_interconnect_0_ram_s1_write,                            --                                   .write
			RAM_s1_read                              => mm_interconnect_0_ram_s1_read,                             --                                   .read
			RAM_s1_readdata                          => mm_interconnect_0_ram_s1_readdata,                         --                                   .readdata
			RAM_s1_writedata                         => mm_interconnect_0_ram_s1_writedata,                        --                                   .writedata
			RAM_s1_byteenable                        => mm_interconnect_0_ram_s1_byteenable,                       --                                   .byteenable
			RAM_s1_readdatavalid                     => mm_interconnect_0_ram_s1_readdatavalid,                    --                                   .readdatavalid
			RAM_s1_waitrequest                       => mm_interconnect_0_ram_s1_waitrequest,                      --                                   .waitrequest
			RAM_s1_chipselect                        => mm_interconnect_0_ram_s1_chipselect,                       --                                   .chipselect
			SPI_MASTER_spi_control_port_address      => mm_interconnect_0_spi_master_spi_control_port_address,     --        SPI_MASTER_spi_control_port.address
			SPI_MASTER_spi_control_port_write        => mm_interconnect_0_spi_master_spi_control_port_write,       --                                   .write
			SPI_MASTER_spi_control_port_read         => mm_interconnect_0_spi_master_spi_control_port_read,        --                                   .read
			SPI_MASTER_spi_control_port_readdata     => mm_interconnect_0_spi_master_spi_control_port_readdata,    --                                   .readdata
			SPI_MASTER_spi_control_port_writedata    => mm_interconnect_0_spi_master_spi_control_port_writedata,   --                                   .writedata
			SPI_MASTER_spi_control_port_chipselect   => mm_interconnect_0_spi_master_spi_control_port_chipselect,  --                                   .chipselect
			SYS_TIMER_s1_address                     => mm_interconnect_0_sys_timer_s1_address,                    --                       SYS_TIMER_s1.address
			SYS_TIMER_s1_write                       => mm_interconnect_0_sys_timer_s1_write,                      --                                   .write
			SYS_TIMER_s1_readdata                    => mm_interconnect_0_sys_timer_s1_readdata,                   --                                   .readdata
			SYS_TIMER_s1_writedata                   => mm_interconnect_0_sys_timer_s1_writedata,                  --                                   .writedata
			SYS_TIMER_s1_chipselect                  => mm_interconnect_0_sys_timer_s1_chipselect,                 --                                   .chipselect
			SYSID_control_slave_address              => mm_interconnect_0_sysid_control_slave_address,             --                SYSID_control_slave.address
			SYSID_control_slave_readdata             => mm_interconnect_0_sysid_control_slave_readdata,            --                                   .readdata
			TS_TIMER_s1_address                      => mm_interconnect_0_ts_timer_s1_address,                     --                        TS_TIMER_s1.address
			TS_TIMER_s1_write                        => mm_interconnect_0_ts_timer_s1_write,                       --                                   .write
			TS_TIMER_s1_readdata                     => mm_interconnect_0_ts_timer_s1_readdata,                    --                                   .readdata
			TS_TIMER_s1_writedata                    => mm_interconnect_0_ts_timer_s1_writedata,                   --                                   .writedata
			TS_TIMER_s1_chipselect                   => mm_interconnect_0_ts_timer_s1_chipselect                   --                                   .chipselect
		);

	irq_mapper : component qsys_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => niosii_irq_irq                  --    sender.irq
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_ram_s1_read_ports_inv <= not mm_interconnect_0_ram_s1_read;

	mm_interconnect_0_ram_s1_byteenable_ports_inv <= not mm_interconnect_0_ram_s1_byteenable;

	mm_interconnect_0_ram_s1_write_ports_inv <= not mm_interconnect_0_ram_s1_write;

	mm_interconnect_0_pio_led_s1_write_ports_inv <= not mm_interconnect_0_pio_led_s1_write;

	mm_interconnect_0_pio_btn_s1_write_ports_inv <= not mm_interconnect_0_pio_btn_s1_write;

	mm_interconnect_0_sys_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_timer_s1_write;

	mm_interconnect_0_ts_timer_s1_write_ports_inv <= not mm_interconnect_0_ts_timer_s1_write;

	mm_interconnect_0_pio_d7seg_s1_write_ports_inv <= not mm_interconnect_0_pio_d7seg_s1_write;

	mm_interconnect_0_spi_master_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_master_spi_control_port_read;

	mm_interconnect_0_spi_master_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_master_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of qsys
